library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity LED_FADING_BLOCK is
    port (
        ck      	: in std_logic;
        reset   	: in std_logic;
        en_led 		: in std_logic;

        color		: out std_logic_vector (23 downto 0);
		en_next_led	: out std_logic
    );
end LED_FADING_BLOCK;

architecture Behavioral of LED_FADING_BLOCK is

	-- Frequency divisor 
	signal cnt_div  													: unsigned (17 downto 0);
	signal ck_en 														: std_logic;
	-- Operations flip -> add/odd -> flip registers
	signal blue_aux, red_aux, green_aux 								: unsigned (7 downto 0);
	signal blue, red, green 											: unsigned (7 downto 0);
	
	-- "Fade color" Finite State machine
	signal en_count_blue, en_count_red, en_count_green					: std_logic;
	signal inc, dec														: std_logic;
	type estado1 is (IDLE1, INC0, INC1, DEC0, INC2, DEC1, INC3, DEC2);
		signal state1, state1_nxt : estado1;
    -- decoder

begin

--- FREQUENCY DIVISOR -----
FREQ_DIV : process (ck, reset)	-- this process outputs ck_en to drive changing of brightness of the chose color
	begin
		if (reset = '1') then
				
			cnt_div <= (others => '0');
			ck_en <= '0';
		
		elsif (ck'event and ck = '1') then
			if (cnt_div < 124999) then		-- IF CHANGED, CHANGE cnt_div AS WELL
				cnt_div <= cnt_div + 1;		-- The frequency for the LED must be > 400 Hz
				ck_en <= '0';
					
			else
				cnt_div <= (others => '0');
				ck_en <= '1';				-- When ck_en = '1', LED assume the current color
			end if;
		end if;
end process;
			

----- FADING AUX  ------  -- flip and add/odd an offset to the color chose by the sequence of the FSM
FLIP_ADD_ODD_AUX : process (ck, reset) 
begin
	if (reset = '1') then
		green_aux 		<= (others => '0');
		red_aux 		<= (others => '0');
		blue_aux 		<= (others => '0');
	elsif (ck'event and ck = '1') then
		if (ck_en = '1') then
			if (en_count_blue = '1') then		-- en_count_blue is generated by the FSM and selects what 8 bit's group must change
				if (inc = '1') then			
					blue_aux <=         		-- Put in an auxiliar signal the sum of blue flipped,
								(blue(0) &		--
								blue(1) &		--
								blue(2) &		--
								blue(3) &		--
								blue(4) &		--
								blue(5) &		--
								blue(6) &		--
								blue(7)) + 5 ;	-- plus an offset (to change the brightness)
				elsif (dec = '1') then
					blue_aux <= 
								(blue(0) &
								blue(1) &
								blue(2) &
								blue(3) &
								blue(4) & 
								blue(5) & 
								blue(6) &
								blue(7)) - 5 ;
				end if;
			elsif (en_count_red = '1') then
				if (inc = '1') then	
					red_aux <= 
								(red(0) &
								red(1) &
								red(2) &
								red(3) &
								red(4) &
								red(5) &
								red(6) &
								red(7)) + 5 ;
				elsif (dec = '1') then
					red_aux <= 
								(red(0) &
								red(1) &
								red(2) &
								red(3) &
								red(4) & 
								red(5) & 
								red(6) &
								red(7)) - 5 ;
				end if;
			elsif (en_count_green = '1') then
				if (inc = '1') then	
					green_aux <= 
								(green(0) &
								green(1) &
								green(2) &
								green(3) &
								green(4) &
								green(5) &
								green(6) &
								green(7)) + 5 ;
				elsif (dec = '1') then
					green_aux <= 
								(green(0) &
								green(1) &
								green(2) &
								green(3) &
								green(4) & 
								green(5) & 
								green(6) &
								green(7)) - 5 ;
				end if;
			end if;
		end if;
	end if;						

end process;
		
------ FADING -----					-- this with the previous process complete the "flip -> add/odd -> flip" function
FLIP_ADD_ODD : process (ck, reset)	-- I want to realize. In particular, this process gets the final reverse operation 
	begin							-- and outputs the color signal.	
		if (reset = '1') then					-- This operation is necessary to respect
			color 	<= (others => '0');			-- the correct order of the bits to send to the LED.
			green 	<= (others => '0');			-- G R B = 7654321_7654321_7654321 where the
			red 	<= (others => '0');			-- rightmost bit of each 8 bit (of each color)
			blue 	<= (others => '0');			-- drive the highest brightness, the leftmost 
		elsif (ck'event and ck = '1') then		-- the lowest one.
			blue 			
					<= blue_aux(0) &
						blue_aux(1) & 
						blue_aux(2) & 
						blue_aux(3) & 
						blue_aux(4) & 
						blue_aux(5) & 
						blue_aux(6) & 
						blue_aux(7);  
			red 			
					<= red_aux(0) &
						red_aux(1) & 
						red_aux(2) & 
						red_aux(3) & 
						red_aux(4) & 
						red_aux(5) & 
						red_aux(6) & 
						red_aux(7);
			green			
					<= green_aux(0) &
						green_aux(1) & 
						green_aux(2) & 
						green_aux(3) & 
						green_aux(4) & 
						green_aux(5) & 
						green_aux(6) & 
						green_aux(7);
		end if;							
		color <= std_logic_vector(blue & red & green);  -- color [23:0] signal
end process;


	

	
	----- FIRST Finite State Machine to control LED fading
	
FADE_LED_FSM : process (ck, reset)  			-- In this FSM I set up a precise sequence to color the LED.
	begin										-- I add and odd bit to reach this sequence:
		if (reset = '1') then					-- 000000->FF0000->FF00FF->0000FF->00FF00->FFFF00->FF0000->...
			state1 <= IDLE1;
		elsif (ck'event and ck = '1') then
			state1 <= state1_nxt;
		end if;
end process;
						
process (blue, red, green, state1, en_led, en_led)
	begin
		case state1 is
			when IDLE1 =>
				if (en_led = '1') then		-- the OR operator is useful to control the
					state1_nxt <= INC0;		-- first LED starting fading and the others.
				else						-- Specifically, "en_led" control the first, 
					state1_nxt <= IDLE1;	-- "en_next_led" control the others for a
				end if;						-- fading sequence
			when INC0 =>					-- starts from state1 = x"000000"
				if (green = "11111111") then
					state1_nxt <= INC1;
				else
					state1_nxt <= INC0;
				end if;
			when INC1 =>					-- starts from state1 = x"FF0000"
				if (blue = "11111111") then
					state1_nxt <= DEC0;
				else
					state1_nxt <= INC1;
				end if;
			when DEC0 =>					-- starts from state1 = x"FF00FF"
				if (green = "00000000") then
					state1_nxt <= INC2;
				else
					state1_nxt <= DEC0;
				end if;
			when INC2 =>					-- starts from state1 = x"0000FF"
				if (red = "11111111") then
					state1_nxt <= DEC1;
				else
					state1_nxt <= INC2; 
				end if;
			when DEC1 =>					-- starts from state1 = x"00FFFF"
				if (blue = "00000000") then
					state1_nxt <= INC3;
				else
					state1_nxt <= DEC1;
				end if;
			when INC3 =>					-- starts from state1 = x"00FF00"
				if (green = "11111111") then
					state1_nxt <= DEC2;
				else
					state1_nxt <= INC3;
				end if;
			when DEC2 =>					-- starts from state1 = x"FFFF00"
				if (red = "00000000") then
					state1_nxt <= INC1;  -- INC1, not INC0 to avoid stepping up a clock cycle
				else
					state1_nxt <= DEC2;  
				end if;
								
			when others => 
				state1_nxt <= IDLE1;
		end case;
end process;
								
process (state1)
	begin
		case state1 is
			when IDLE1 =>            
					inc       			<= '0';	-- A possible future implementation can be to make a control here
					dec       			<= '0';	-- on the "color" signal of the top level module to allow,
					en_count_blue 		<= '0';	-- when I click the button to change the fading mode, that
					en_count_red 		<= '0';	-- this one starts over from the last "color" value. It can
					en_count_green 		<= '0';	-- be implemented by a if-else construct that brigngs you
					en_next_led 		<= '0';	-- directly to the right color in the states
			when INC0 =>				
					inc       			<= '1';
					dec       			<= '0';
					en_count_blue 		<= '0';
					en_count_red 		<= '0';
					en_count_green 		<= '1';
					if (green = "11111111") then
						en_next_led <= '1';	-- I want this sequence: when the current LED is "FF0000",
					else					-- the previous LED will be at "000000",
						en_next_led <= '0';	-- and the next LED of the current one is "FF00FF"
					end if; 
			when INC1 =>				
					inc       			<= '1';
					dec       			<= '0';
					en_count_blue 		<= '1';
					en_count_red 		<= '0';
					en_count_green 		<= '0';
					en_next_led 		<= '0';
			when DEC0 =>				
					inc       			<= '0';
					dec       			<= '1';
					en_count_blue 		<= '0';
					en_count_red 		<= '0';
					en_count_green 		<= '1';
					en_next_led 		<= '0';
			when INC2 =>				
					inc       			<= '1';
					dec       			<= '0';
					en_count_blue 		<= '0';
					en_count_red 		<= '1';
					en_count_green 		<= '0';
					en_next_led 		<= '0';
			when DEC1 =>				
					inc       			<= '0';
					dec       			<= '1';
					en_count_blue 		<= '1';
					en_count_red 		<= '0';
					en_count_green 		<= '0';
					en_next_led 		<= '0';
			when INC3 =>				
					inc       			<= '1';
					dec       			<= '0';
					en_count_blue 		<= '0';
					en_count_red 		<= '0';
					en_count_green 		<= '1';
					en_next_led 		<= '0';
			when DEC2 =>				
					inc       			<= '0';
					dec       			<= '1';
					en_count_blue 		<= '0';
					en_count_red 		<= '1';
					en_count_green 		<= '0';
					en_next_led 		<= '0';
				 
			when others => 
					inc       			<= '0';
					dec       			<= '0';
					en_count_blue 		<= '0';
					en_count_red 		<= '0';
					en_count_green 		<= '0';
					en_next_led 		<= '0';
		end case;
end process;

end Behavioral;